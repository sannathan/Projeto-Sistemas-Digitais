module seletor(a, b, sinal_a, sinal_b, botao_1, botao_2, botao_3, botao_4, clk, saida, sinal_saida);